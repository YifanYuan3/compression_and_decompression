`define DATA_WIDTH 256

module Compressor (
	input [DATA_WIDTH - 1: 0] data;
);


endmodule